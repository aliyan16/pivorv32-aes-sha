

module Inv_mix_cols(output [127:0] Dout, input [127:0] Din);


	wire [7:0] b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15;
	reg [7:0] S3, S2, S1, S0, C0, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15;

	assign b0 = Din[7:0];
	assign b1 = Din[15:8];
	assign b2 = Din[23:16];
	assign b3 = Din[31:24];
	assign b4 = Din[39:32];
	assign b5 = Din[47:40];
	assign b6 = Din[55:48];
	assign b7 = Din[63:56];
	assign b8 = Din[71:64];
	assign b9 = Din[79:72];
	assign b10 = Din[87:80];
	assign b11 = Din[95:88];
	assign b12 = Din[103:96];
	assign b13 = Din[111:104];
	assign b14 = Din[119:112];
	assign b15 = Din[127:120];
	
	assign Dout[7:0] = C0;
	assign Dout[15:8] = C1;
	assign Dout[23:16] = C2;
	assign Dout[31:24] = C3;
	assign Dout[39:32] = C4;
	assign Dout[47:40] = C5;
	assign Dout[55:48] = C6;
	assign Dout[63:56] = C7;
	assign Dout[71:64] = C8;
	assign Dout[79:72] = C9;
	assign Dout[87:80] = C10;
	assign Dout[95:88] = C11;
	assign Dout[103:96] = C12;
	assign Dout[111:104] = C13;
	assign Dout[119:112] = C14;
	assign Dout[127:120] = C15;
	
	
	always @(*) begin
		S3 = multiply(b15, 14);
		S2 = multiply(b14, 11);
		S1 = multiply(b13, 13);
		S0 = multiply(b12, 9);
		C15 = multiply(b15, 14) ^ multiply(b14, 11) ^ multiply(b13, 13) ^ multiply(b12, 9);
		C14 = multiply(b15, 9) ^ multiply(b14, 14) ^ multiply(b13, 11) ^ multiply(b12, 13);
		C13 = multiply(b15, 13) ^ multiply(b14, 9) ^ multiply(b13, 14) ^ multiply(b12, 11);
		C12 = multiply(b15, 11) ^ multiply(b14, 13) ^ multiply(b13, 9) ^ multiply(b12, 14);		

		C11 = multiply(b11, 14) ^ multiply(b10, 11) ^ multiply(b9, 13) ^ multiply(b8, 9);
		C10 = multiply(b11, 9) ^ multiply(b10, 14) ^ multiply(b9, 11) ^ multiply(b8, 13);
		C9 = multiply(b11, 13) ^ multiply(b10, 9) ^ multiply(b9, 14) ^ multiply(b8, 11);
		C8 = multiply(b11, 11) ^ multiply(b10, 13) ^ multiply(b9, 9) ^ multiply(b8, 14);

		C7 = multiply(b7, 14) ^ multiply(b6, 11) ^ multiply(b5, 13) ^ multiply(b4, 9);
		C6 = multiply(b7, 9) ^ multiply(b6, 14) ^ multiply(b5, 11) ^ multiply(b4, 13);
		C5 = multiply(b7, 13) ^ multiply(b6, 9) ^ multiply(b5, 14) ^ multiply(b4, 11);
		C4 = multiply(b7, 11) ^ multiply(b6, 13) ^ multiply(b5, 9) ^ multiply(b4, 14);

		C3 = multiply(b3, 14) ^ multiply(b2, 11) ^ multiply(b1, 13) ^ multiply(b0, 9);
		C2 = multiply(b3, 9) ^ multiply(b2, 14) ^ multiply(b1, 11) ^ multiply(b0, 13);
		C1 = multiply(b3, 13) ^ multiply(b2, 9) ^ multiply(b1, 14) ^ multiply(b0, 11);
		C0 = multiply(b3, 11) ^ multiply(b2, 13) ^ multiply(b1, 9) ^ multiply(b0, 14);
	end
	
	function integer multiply (input integer a, input integer b);
			if (b == 9)
				multiply = lut_9(a);
			else if (b == 11)
				multiply = lut_11(a);
			else if (b == 13)
				multiply = lut_13(a);
			else if (b == 14)
				multiply = lut_14(a);
	endfunction
	
	function integer lut_9(input integer a);
		case (a)
			8'h00: lut_9 = 8'h00;
			8'h01: lut_9 = 8'h09;
			8'h02: lut_9 = 8'h12;
			8'h03: lut_9 = 8'h1B;
			8'h04: lut_9 = 8'h24;
			8'h05: lut_9 = 8'h2D;
			8'h06: lut_9 = 8'h36;
			8'h07: lut_9 = 8'h3F;
			8'h08: lut_9 = 8'h48;
			8'h09: lut_9 = 8'h41;
			8'h0A: lut_9 = 8'h5A;
			8'h0B: lut_9 = 8'h53;
			8'h0C: lut_9 = 8'h6C;
			8'h0D: lut_9 = 8'h65;
			8'h0E: lut_9 = 8'h7E;
			8'h0F: lut_9 = 8'h77;
			8'h10: lut_9 = 8'h90;
			8'h11: lut_9 = 8'h99;
			8'h12: lut_9 = 8'h82;
			8'h13: lut_9 = 8'h8B;
			8'h14: lut_9 = 8'hB4;
			8'h15: lut_9 = 8'hBD;
			8'h16: lut_9 = 8'hA6;
			8'h17: lut_9 = 8'hAF;
			8'h18: lut_9 = 8'hD8;
			8'h19: lut_9 = 8'hD1;
			8'h1A: lut_9 = 8'hCA;
			8'h1B: lut_9 = 8'hC3;
			8'h1C: lut_9 = 8'hFC;
			8'h1D: lut_9 = 8'hF5;
			8'h1E: lut_9 = 8'hEE;
			8'h1F: lut_9 = 8'hE7;
			8'h20: lut_9 = 8'h3B;
			8'h21: lut_9 = 8'h32;
			8'h22: lut_9 = 8'h29;
			8'h23: lut_9 = 8'h20;
			8'h24: lut_9 = 8'h1F;
			8'h25: lut_9 = 8'h16;
			8'h26: lut_9 = 8'h0D;
			8'h27: lut_9 = 8'h04;
			8'h28: lut_9 = 8'h73;
			8'h29: lut_9 = 8'h7A;
			8'h2A: lut_9 = 8'h61;
			8'h2B: lut_9 = 8'h68;
			8'h2C: lut_9 = 8'h57;
			8'h2D: lut_9 = 8'h5E;
			8'h2E: lut_9 = 8'h45;
			8'h2F: lut_9 = 8'h4C;
			8'h30: lut_9 = 8'hAB;
			8'h31: lut_9 = 8'hA2;
			8'h32: lut_9 = 8'hB9;
			8'h33: lut_9 = 8'hB0;
			8'h34: lut_9 = 8'h8F;
			8'h35: lut_9 = 8'h86;
			8'h36: lut_9 = 8'h9D;
			8'h37: lut_9 = 8'h94;
			8'h38: lut_9 = 8'hE3;
			8'h39: lut_9 = 8'hEA;
			8'h3A: lut_9 = 8'hF1;
			8'h3B: lut_9 = 8'hF8;
			8'h3C: lut_9 = 8'hC7;
			8'h3D: lut_9 = 8'hCE;
			8'h3E: lut_9 = 8'hD5;
			8'h3F: lut_9 = 8'hDC;
			8'h40: lut_9 = 8'h76;
			8'h41: lut_9 = 8'h7F;
			8'h42: lut_9 = 8'h64;
			8'h43: lut_9 = 8'h6D;
			8'h44: lut_9 = 8'h52;
			8'h45: lut_9 = 8'h5B;
			8'h46: lut_9 = 8'h40;
			8'h47: lut_9 = 8'h49;
			8'h48: lut_9 = 8'h3E;
			8'h49: lut_9 = 8'h37;
			8'h4A: lut_9 = 8'h2C;
			8'h4B: lut_9 = 8'h25;
			8'h4C: lut_9 = 8'h1A;
			8'h4D: lut_9 = 8'h13;
			8'h4E: lut_9 = 8'h08;
			8'h4F: lut_9 = 8'h01;
			8'h50: lut_9 = 8'hE6;
			8'h51: lut_9 = 8'hEF;
			8'h52: lut_9 = 8'hF4;
			8'h53: lut_9 = 8'hFD;
			8'h54: lut_9 = 8'hC2;
			8'h55: lut_9 = 8'hCB;
			8'h56: lut_9 = 8'hD0;
			8'h57: lut_9 = 8'hD9;
			8'h58: lut_9 = 8'hAE;
			8'h59: lut_9 = 8'hA7;
			8'h5A: lut_9 = 8'hBC;
			8'h5B: lut_9 = 8'hB5;
			8'h5C: lut_9 = 8'h8A;
			8'h5D: lut_9 = 8'h83;
			8'h5E: lut_9 = 8'h98;
			8'h5F: lut_9 = 8'h91;
			8'h60: lut_9 = 8'h4D;
			8'h61: lut_9 = 8'h44;
			8'h62: lut_9 = 8'h5F;
			8'h63: lut_9 = 8'h56;
			8'h64: lut_9 = 8'h69;
			8'h65: lut_9 = 8'h60;
			8'h66: lut_9 = 8'h7B;
			8'h67: lut_9 = 8'h72;
			8'h68: lut_9 = 8'h05;
			8'h69: lut_9 = 8'h0C;
			8'h6A: lut_9 = 8'h17;
			8'h6B: lut_9 = 8'h1E;
			8'h6C: lut_9 = 8'h21;
			8'h6D: lut_9 = 8'h28;
			8'h6E: lut_9 = 8'h33;
			8'h6F: lut_9 = 8'h3A;
			8'h70: lut_9 = 8'hDD;
			8'h71: lut_9 = 8'hD4;
			8'h72: lut_9 = 8'hCF;
			8'h73: lut_9 = 8'hC6;
			8'h74: lut_9 = 8'hF9;
			8'h75: lut_9 = 8'hF0;
			8'h76: lut_9 = 8'hEB;
			8'h77: lut_9 = 8'hE2;
			8'h78: lut_9 = 8'h95;
			8'h79: lut_9 = 8'h9C;
			8'h7A: lut_9 = 8'h87;
			8'h7B: lut_9 = 8'h8E;
			8'h7C: lut_9 = 8'hB1;
			8'h7D: lut_9 = 8'hB8;
			8'h7E: lut_9 = 8'hA3;
			8'h7F: lut_9 = 8'hAA;
			8'h80: lut_9 = 8'hEC;
			8'h81: lut_9 = 8'hE5;
			8'h82: lut_9 = 8'hFE;
			8'h83: lut_9 = 8'hF7;
			8'h84: lut_9 = 8'hC8;
			8'h85: lut_9 = 8'hC1;
			8'h86: lut_9 = 8'hDA;
			8'h87: lut_9 = 8'hD3;
			8'h88: lut_9 = 8'hA4;
			8'h89: lut_9 = 8'hAD;
			8'h8A: lut_9 = 8'hB6;
			8'h8B: lut_9 = 8'hBF;
			8'h8C: lut_9 = 8'h80;
			8'h8D: lut_9 = 8'h89;
			8'h8E: lut_9 = 8'h92;
			8'h8F: lut_9 = 8'h9B;
			8'h90: lut_9 = 8'h7C;
			8'h91: lut_9 = 8'h75;
			8'h92: lut_9 = 8'h6E;
			8'h93: lut_9 = 8'h67;
			8'h94: lut_9 = 8'h58;
			8'h95: lut_9 = 8'h51;
			8'h96: lut_9 = 8'h4A;
			8'h97: lut_9 = 8'h43;
			8'h98: lut_9 = 8'h34;
			8'h99: lut_9 = 8'h3D;
			8'h9A: lut_9 = 8'h26;
			8'h9B: lut_9 = 8'h2F;
			8'h9C: lut_9 = 8'h10;
			8'h9D: lut_9 = 8'h19;
			8'h9E: lut_9 = 8'h02;
			8'h9F: lut_9 = 8'h0B;
			8'hA0: lut_9 = 8'hD7;
			8'hA1: lut_9 = 8'hDE;
			8'hA2: lut_9 = 8'hC5;
			8'hA3: lut_9 = 8'hCC;
			8'hA4: lut_9 = 8'hF3;
			8'hA5: lut_9 = 8'hFA;
			8'hA6: lut_9 = 8'hE1;
			8'hA7: lut_9 = 8'hE8;
			8'hA8: lut_9 = 8'h9F;
			8'hA9: lut_9 = 8'h96;
			8'hAA: lut_9 = 8'h8D;
			8'hAB: lut_9 = 8'h84;
			8'hAC: lut_9 = 8'hBB;
			8'hAD: lut_9 = 8'hB2;
			8'hAE: lut_9 = 8'hA9;
			8'hAF: lut_9 = 8'hA0;
			8'hB0: lut_9 = 8'h47;
			8'hB1: lut_9 = 8'h4E;
			8'hB2: lut_9 = 8'h55;
			8'hB3: lut_9 = 8'h5C;
			8'hB4: lut_9 = 8'h63;
			8'hB5: lut_9 = 8'h6A;
			8'hB6: lut_9 = 8'h71;
			8'hB7: lut_9 = 8'h78;
			8'hB8: lut_9 = 8'h0F;
			8'hB9: lut_9 = 8'h06;
			8'hBA: lut_9 = 8'h1D;
			8'hBB: lut_9 = 8'h14;
			8'hBC: lut_9 = 8'h2B;
			8'hBD: lut_9 = 8'h22;
			8'hBE: lut_9 = 8'h39;
			8'hBF: lut_9 = 8'h30;
			8'hC0: lut_9 = 8'h9A;
			8'hC1: lut_9 = 8'h93;
			8'hC2: lut_9 = 8'h88;
			8'hC3: lut_9 = 8'h81;
			8'hC4: lut_9 = 8'hBE;
			8'hC5: lut_9 = 8'hB7;
			8'hC6: lut_9 = 8'hAC;
			8'hC7: lut_9 = 8'hA5;
			8'hC8: lut_9 = 8'hD2;
			8'hC9: lut_9 = 8'hDB;
			8'hCA: lut_9 = 8'hC0;
			8'hCB: lut_9 = 8'hC9;
			8'hCC: lut_9 = 8'hF6;
			8'hCD: lut_9 = 8'hFF;
			8'hCE: lut_9 = 8'hE4;
			8'hCF: lut_9 = 8'hED;
			8'hD0: lut_9 = 8'h0A;
			8'hD1: lut_9 = 8'h03;
			8'hD2: lut_9 = 8'h18;
			8'hD3: lut_9 = 8'h11;
			8'hD4: lut_9 = 8'h2E;
			8'hD5: lut_9 = 8'h27;
			8'hD6: lut_9 = 8'h3C;
			8'hD7: lut_9 = 8'h35;
			8'hD8: lut_9 = 8'h42;
			8'hD9: lut_9 = 8'h4B;
			8'hDA: lut_9 = 8'h50;
			8'hDB: lut_9 = 8'h59;
			8'hDC: lut_9 = 8'h66;
			8'hDD: lut_9 = 8'h6F;
			8'hDE: lut_9 = 8'h74;
			8'hDF: lut_9 = 8'h7D;
			8'hE0: lut_9 = 8'hA1;
			8'hE1: lut_9 = 8'hA8;
			8'hE2: lut_9 = 8'hB3;
			8'hE3: lut_9 = 8'hBA;
			8'hE4: lut_9 = 8'h85;
			8'hE5: lut_9 = 8'h8C;
			8'hE6: lut_9 = 8'h97;
			8'hE7: lut_9 = 8'h9E;
			8'hE8: lut_9 = 8'hE9;
			8'hE9: lut_9 = 8'hE0;
			8'hEA: lut_9 = 8'hFB;
			8'hEB: lut_9 = 8'hF2;
			8'hEC: lut_9 = 8'hCD;
			8'hED: lut_9 = 8'hC4;
			8'hEE: lut_9 = 8'hDF;
			8'hEF: lut_9 = 8'hD6;
			8'hF0: lut_9 = 8'h31;
			8'hF1: lut_9 = 8'h38;
			8'hF2: lut_9 = 8'h23;
			8'hF3: lut_9 = 8'h2A;
			8'hF4: lut_9 = 8'h15;
			8'hF5: lut_9 = 8'h1C;
			8'hF6: lut_9 = 8'h07;
			8'hF7: lut_9 = 8'h0E;
			8'hF8: lut_9 = 8'h79;
			8'hF9: lut_9 = 8'h70;
			8'hFA: lut_9 = 8'h6B;
			8'hFB: lut_9 = 8'h62;
			8'hFC: lut_9 = 8'h5D;
			8'hFD: lut_9 = 8'h54;
			8'hFE: lut_9 = 8'h4F;
			default: lut_9 = 8'h46;
		endcase
	endfunction
	
	function integer lut_11(input integer a);
		case (a)
			8'h00: lut_11 = 8'h00;
			8'h01: lut_11 = 8'h0B;
			8'h02: lut_11 = 8'h16;
			8'h03: lut_11 = 8'h1D;
			8'h04: lut_11 = 8'h2C;
			8'h05: lut_11 = 8'h27;
			8'h06: lut_11 = 8'h3A;
			8'h07: lut_11 = 8'h31;
			8'h08: lut_11 = 8'h58;
			8'h09: lut_11 = 8'h53;
			8'h0A: lut_11 = 8'h4E;
			8'h0B: lut_11 = 8'h45;
			8'h0C: lut_11 = 8'h74;
			8'h0D: lut_11 = 8'h7F;
			8'h0E: lut_11 = 8'h62;
			8'h0F: lut_11 = 8'h69;
			8'h10: lut_11 = 8'hB0;
			8'h11: lut_11 = 8'hBB;
			8'h12: lut_11 = 8'hA6;
			8'h13: lut_11 = 8'hAD;
			8'h14: lut_11 = 8'h9C;
			8'h15: lut_11 = 8'h97;
			8'h16: lut_11 = 8'h8A;
			8'h17: lut_11 = 8'h81;
			8'h18: lut_11 = 8'hE8;
			8'h19: lut_11 = 8'hE3;
			8'h1A: lut_11 = 8'hFE;
			8'h1B: lut_11 = 8'hF5;
			8'h1C: lut_11 = 8'hC4;
			8'h1D: lut_11 = 8'hCF;
			8'h1E: lut_11 = 8'hD2;
			8'h1F: lut_11 = 8'hD9;
			8'h20: lut_11 = 8'h7B;
			8'h21: lut_11 = 8'h70;
			8'h22: lut_11 = 8'h6D;
			8'h23: lut_11 = 8'h66;
			8'h24: lut_11 = 8'h57;
			8'h25: lut_11 = 8'h5C;
			8'h26: lut_11 = 8'h41;
			8'h27: lut_11 = 8'h4A;
			8'h28: lut_11 = 8'h23;
			8'h29: lut_11 = 8'h28;
			8'h2A: lut_11 = 8'h35;
			8'h2B: lut_11 = 8'h3E;
			8'h2C: lut_11 = 8'h0F;
			8'h2D: lut_11 = 8'h04;
			8'h2E: lut_11 = 8'h19;
			8'h2F: lut_11 = 8'h12;
			8'h30: lut_11 = 8'hCB;
			8'h31: lut_11 = 8'hC0;
			8'h32: lut_11 = 8'hDD;
			8'h33: lut_11 = 8'hD6;
			8'h34: lut_11 = 8'hE7;
			8'h35: lut_11 = 8'hEC;
			8'h36: lut_11 = 8'hF1;
			8'h37: lut_11 = 8'hFA;
			8'h38: lut_11 = 8'h93;
			8'h39: lut_11 = 8'h98;
			8'h3A: lut_11 = 8'h85;
			8'h3B: lut_11 = 8'h8E;
			8'h3C: lut_11 = 8'hBF;
			8'h3D: lut_11 = 8'hB4;
			8'h3E: lut_11 = 8'hA9;
			8'h3F: lut_11 = 8'hA2;
			8'h40: lut_11 = 8'hF6;
			8'h41: lut_11 = 8'hFD;
			8'h42: lut_11 = 8'hE0;
			8'h43: lut_11 = 8'hEB;
			8'h44: lut_11 = 8'hDA;
			8'h45: lut_11 = 8'hD1;
			8'h46: lut_11 = 8'hCC;
			8'h47: lut_11 = 8'hC7;
			8'h48: lut_11 = 8'hAE;
			8'h49: lut_11 = 8'hA5;
			8'h4A: lut_11 = 8'hB8;
			8'h4B: lut_11 = 8'hB3;
			8'h4C: lut_11 = 8'h82;
			8'h4D: lut_11 = 8'h89;
			8'h4E: lut_11 = 8'h94;
			8'h4F: lut_11 = 8'h9F;
			8'h50: lut_11 = 8'h46;
			8'h51: lut_11 = 8'h4D;
			8'h52: lut_11 = 8'h50;
			8'h53: lut_11 = 8'h5B;
			8'h54: lut_11 = 8'h6A;
			8'h55: lut_11 = 8'h61;
			8'h56: lut_11 = 8'h7C;
			8'h57: lut_11 = 8'h77;
			8'h58: lut_11 = 8'h1E;
			8'h59: lut_11 = 8'h15;
			8'h5A: lut_11 = 8'h08;
			8'h5B: lut_11 = 8'h03;
			8'h5C: lut_11 = 8'h32;
			8'h5D: lut_11 = 8'h39;
			8'h5E: lut_11 = 8'h24;
			8'h5F: lut_11 = 8'h2F;
			8'h60: lut_11 = 8'h8D;
			8'h61: lut_11 = 8'h86;
			8'h62: lut_11 = 8'h9B;
			8'h63: lut_11 = 8'h90;
			8'h64: lut_11 = 8'hA1;
			8'h65: lut_11 = 8'hAA;
			8'h66: lut_11 = 8'hB7;
			8'h67: lut_11 = 8'hBC;
			8'h68: lut_11 = 8'hD5;
			8'h69: lut_11 = 8'hDE;
			8'h6A: lut_11 = 8'hC3;
			8'h6B: lut_11 = 8'hC8;
			8'h6C: lut_11 = 8'hF9;
			8'h6D: lut_11 = 8'hF2;
			8'h6E: lut_11 = 8'hEF;
			8'h6F: lut_11 = 8'hE4;
			8'h70: lut_11 = 8'h3D;
			8'h71: lut_11 = 8'h36;
			8'h72: lut_11 = 8'h2B;
			8'h73: lut_11 = 8'h20;
			8'h74: lut_11 = 8'h11;
			8'h75: lut_11 = 8'h1A;
			8'h76: lut_11 = 8'h07;
			8'h77: lut_11 = 8'h0C;
			8'h78: lut_11 = 8'h65;
			8'h79: lut_11 = 8'h6E;
			8'h7A: lut_11 = 8'h73;
			8'h7B: lut_11 = 8'h78;
			8'h7C: lut_11 = 8'h49;
			8'h7D: lut_11 = 8'h42;
			8'h7E: lut_11 = 8'h5F;
			8'h7F: lut_11 = 8'h54;
			8'h80: lut_11 = 8'hF7;
			8'h81: lut_11 = 8'hFC;
			8'h82: lut_11 = 8'hE1;
			8'h83: lut_11 = 8'hEA;
			8'h84: lut_11 = 8'hDB;
			8'h85: lut_11 = 8'hD0;
			8'h86: lut_11 = 8'hCD;
			8'h87: lut_11 = 8'hC6;
			8'h88: lut_11 = 8'hAF;
			8'h89: lut_11 = 8'hA4;
			8'h8A: lut_11 = 8'hB9;
			8'h8B: lut_11 = 8'hB2;
			8'h8C: lut_11 = 8'h83;
			8'h8D: lut_11 = 8'h88;
			8'h8E: lut_11 = 8'h95;
			8'h8F: lut_11 = 8'h9E;
			8'h90: lut_11 = 8'h47;
			8'h91: lut_11 = 8'h4C;
			8'h92: lut_11 = 8'h51;
			8'h93: lut_11 = 8'h5A;
			8'h94: lut_11 = 8'h6B;
			8'h95: lut_11 = 8'h60;
			8'h96: lut_11 = 8'h7D;
			8'h97: lut_11 = 8'h76;
			8'h98: lut_11 = 8'h1F;
			8'h99: lut_11 = 8'h14;
			8'h9A: lut_11 = 8'h09;
			8'h9B: lut_11 = 8'h02;
			8'h9C: lut_11 = 8'h33;
			8'h9D: lut_11 = 8'h38;
			8'h9E: lut_11 = 8'h25;
			8'h9F: lut_11 = 8'h2E;
			8'hA0: lut_11 = 8'h8C;
			8'hA1: lut_11 = 8'h87;
			8'hA2: lut_11 = 8'h9A;
			8'hA3: lut_11 = 8'h91;
			8'hA4: lut_11 = 8'hA0;
			8'hA5: lut_11 = 8'hAB;
			8'hA6: lut_11 = 8'hB6;
			8'hA7: lut_11 = 8'hBD;
			8'hA8: lut_11 = 8'hD4;
			8'hA9: lut_11 = 8'hDF;
			8'hAA: lut_11 = 8'hC2;
			8'hAB: lut_11 = 8'hC9;
			8'hAC: lut_11 = 8'hF8;
			8'hAD: lut_11 = 8'hF3;
			8'hAE: lut_11 = 8'hEE;
			8'hAF: lut_11 = 8'hE5;
			8'hB0: lut_11 = 8'h3C;
			8'hB1: lut_11 = 8'h37;
			8'hB2: lut_11 = 8'h2A;
			8'hB3: lut_11 = 8'h21;
			8'hB4: lut_11 = 8'h10;
			8'hB5: lut_11 = 8'h1B;
			8'hB6: lut_11 = 8'h06;
			8'hB7: lut_11 = 8'h0D;
			8'hB8: lut_11 = 8'h64;
			8'hB9: lut_11 = 8'h6F;
			8'hBA: lut_11 = 8'h72;
			8'hBB: lut_11 = 8'h79;
			8'hBC: lut_11 = 8'h48;
			8'hBD: lut_11 = 8'h43;
			8'hBE: lut_11 = 8'h5E;
			8'hBF: lut_11 = 8'h55;
			8'hC0: lut_11 = 8'h01;
			8'hC1: lut_11 = 8'h0A;
			8'hC2: lut_11 = 8'h17;
			8'hC3: lut_11 = 8'h1C;
			8'hC4: lut_11 = 8'h2D;
			8'hC5: lut_11 = 8'h26;
			8'hC6: lut_11 = 8'h3B;
			8'hC7: lut_11 = 8'h30;
			8'hC8: lut_11 = 8'h59;
			8'hC9: lut_11 = 8'h52;
			8'hCA: lut_11 = 8'h4F;
			8'hCB: lut_11 = 8'h44;
			8'hCC: lut_11 = 8'h75;
			8'hCD: lut_11 = 8'h7E;
			8'hCE: lut_11 = 8'h63;
			8'hCF: lut_11 = 8'h68;
			8'hD0: lut_11 = 8'hB1;
			8'hD1: lut_11 = 8'hBA;
			8'hD2: lut_11 = 8'hA7;
			8'hD3: lut_11 = 8'hAC;
			8'hD4: lut_11 = 8'h9D;
			8'hD5: lut_11 = 8'h96;
			8'hD6: lut_11 = 8'h8B;
			8'hD7: lut_11 = 8'h80;
			8'hD8: lut_11 = 8'hE9;
			8'hD9: lut_11 = 8'hE2;
			8'hDA: lut_11 = 8'hFF;
			8'hDB: lut_11 = 8'hF4;
			8'hDC: lut_11 = 8'hC5;
			8'hDD: lut_11 = 8'hCE;
			8'hDE: lut_11 = 8'hD3;
			8'hDF: lut_11 = 8'hD8;
			8'hE0: lut_11 = 8'h7A;
			8'hE1: lut_11 = 8'h71;
			8'hE2: lut_11 = 8'h6C;
			8'hE3: lut_11 = 8'h67;
			8'hE4: lut_11 = 8'h56;
			8'hE5: lut_11 = 8'h5D;
			8'hE6: lut_11 = 8'h40;
			8'hE7: lut_11 = 8'h4B;
			8'hE8: lut_11 = 8'h22;
			8'hE9: lut_11 = 8'h29;
			8'hEA: lut_11 = 8'h34;
			8'hEB: lut_11 = 8'h3F;
			8'hEC: lut_11 = 8'h0E;
			8'hED: lut_11 = 8'h05;
			8'hEE: lut_11 = 8'h18;
			8'hEF: lut_11 = 8'h13;
			8'hF0: lut_11 = 8'hCA;
			8'hF1: lut_11 = 8'hC1;
			8'hF2: lut_11 = 8'hDC;
			8'hF3: lut_11 = 8'hD7;
			8'hF4: lut_11 = 8'hE6;
			8'hF5: lut_11 = 8'hED;
			8'hF6: lut_11 = 8'hF0;
			8'hF7: lut_11 = 8'hFB;
			8'hF8: lut_11 = 8'h92;
			8'hF9: lut_11 = 8'h99;
			8'hFA: lut_11 = 8'h84;
			8'hFB: lut_11 = 8'h8F;
			8'hFC: lut_11 = 8'hBE;
			8'hFD: lut_11 = 8'hB5;
			8'hFE: lut_11 = 8'hA8;
			default: lut_11 = 8'hA3;
		endcase
	endfunction
	
	function integer lut_13(input integer a);
		case (a)
			8'h00: lut_13 = 8'h00;
			8'h01: lut_13 = 8'h0D;
			8'h02: lut_13 = 8'h1A;
			8'h03: lut_13 = 8'h17;
			8'h04: lut_13 = 8'h34;
			8'h05: lut_13 = 8'h39;
			8'h06: lut_13 = 8'h2E;
			8'h07: lut_13 = 8'h23;
			8'h08: lut_13 = 8'h68;
			8'h09: lut_13 = 8'h65;
			8'h0A: lut_13 = 8'h72;
			8'h0B: lut_13 = 8'h7F;
			8'h0C: lut_13 = 8'h5C;
			8'h0D: lut_13 = 8'h51;
			8'h0E: lut_13 = 8'h46;
			8'h0F: lut_13 = 8'h4B;
			8'h10: lut_13 = 8'hD0;
			8'h11: lut_13 = 8'hDD;
			8'h12: lut_13 = 8'hCA;
			8'h13: lut_13 = 8'hC7;
			8'h14: lut_13 = 8'hE4;
			8'h15: lut_13 = 8'hE9;
			8'h16: lut_13 = 8'hFE;
			8'h17: lut_13 = 8'hF3;
			8'h18: lut_13 = 8'hB8;
			8'h19: lut_13 = 8'hB5;
			8'h1A: lut_13 = 8'hA2;
			8'h1B: lut_13 = 8'hAF;
			8'h1C: lut_13 = 8'h8C;
			8'h1D: lut_13 = 8'h81;
			8'h1E: lut_13 = 8'h96;
			8'h1F: lut_13 = 8'h9B;
			8'h20: lut_13 = 8'hBB;
			8'h21: lut_13 = 8'hB6;
			8'h22: lut_13 = 8'hA1;
			8'h23: lut_13 = 8'hAC;
			8'h24: lut_13 = 8'h8F;
			8'h25: lut_13 = 8'h82;
			8'h26: lut_13 = 8'h95;
			8'h27: lut_13 = 8'h98;
			8'h28: lut_13 = 8'hD3;
			8'h29: lut_13 = 8'hDE;
			8'h2A: lut_13 = 8'hC9;
			8'h2B: lut_13 = 8'hC4;
			8'h2C: lut_13 = 8'hE7;
			8'h2D: lut_13 = 8'hEA;
			8'h2E: lut_13 = 8'hFD;
			8'h2F: lut_13 = 8'hF0;
			8'h30: lut_13 = 8'h6B;
			8'h31: lut_13 = 8'h66;
			8'h32: lut_13 = 8'h71;
			8'h33: lut_13 = 8'h7C;
			8'h34: lut_13 = 8'h5F;
			8'h35: lut_13 = 8'h52;
			8'h36: lut_13 = 8'h45;
			8'h37: lut_13 = 8'h48;
			8'h38: lut_13 = 8'h03;
			8'h39: lut_13 = 8'h0E;
			8'h3A: lut_13 = 8'h19;
			8'h3B: lut_13 = 8'h14;
			8'h3C: lut_13 = 8'h37;
			8'h3D: lut_13 = 8'h3A;
			8'h3E: lut_13 = 8'h2D;
			8'h3F: lut_13 = 8'h20;
			8'h40: lut_13 = 8'h6D;
			8'h41: lut_13 = 8'h60;
			8'h42: lut_13 = 8'h77;
			8'h43: lut_13 = 8'h7A;
			8'h44: lut_13 = 8'h59;
			8'h45: lut_13 = 8'h54;
			8'h46: lut_13 = 8'h43;
			8'h47: lut_13 = 8'h4E;
			8'h48: lut_13 = 8'h05;
			8'h49: lut_13 = 8'h08;
			8'h4A: lut_13 = 8'h1F;
			8'h4B: lut_13 = 8'h12;
			8'h4C: lut_13 = 8'h31;
			8'h4D: lut_13 = 8'h3C;
			8'h4E: lut_13 = 8'h2B;
			8'h4F: lut_13 = 8'h26;
			8'h50: lut_13 = 8'hBD;
			8'h51: lut_13 = 8'hB0;
			8'h52: lut_13 = 8'hA7;
			8'h53: lut_13 = 8'hAA;
			8'h54: lut_13 = 8'h89;
			8'h55: lut_13 = 8'h84;
			8'h56: lut_13 = 8'h93;
			8'h57: lut_13 = 8'h9E;
			8'h58: lut_13 = 8'hD5;
			8'h59: lut_13 = 8'hD8;
			8'h5A: lut_13 = 8'hCF;
			8'h5B: lut_13 = 8'hC2;
			8'h5C: lut_13 = 8'hE1;
			8'h5D: lut_13 = 8'hEC;
			8'h5E: lut_13 = 8'hFB;
			8'h5F: lut_13 = 8'hF6;
			8'h60: lut_13 = 8'hD6;
			8'h61: lut_13 = 8'hDB;
			8'h62: lut_13 = 8'hCC;
			8'h63: lut_13 = 8'hC1;
			8'h64: lut_13 = 8'hE2;
			8'h65: lut_13 = 8'hEF;
			8'h66: lut_13 = 8'hF8;
			8'h67: lut_13 = 8'hF5;
			8'h68: lut_13 = 8'hBE;
			8'h69: lut_13 = 8'hB3;
			8'h6A: lut_13 = 8'hA4;
			8'h6B: lut_13 = 8'hA9;
			8'h6C: lut_13 = 8'h8A;
			8'h6D: lut_13 = 8'h87;
			8'h6E: lut_13 = 8'h90;
			8'h6F: lut_13 = 8'h9D;
			8'h70: lut_13 = 8'h06;
			8'h71: lut_13 = 8'h0B;
			8'h72: lut_13 = 8'h1C;
			8'h73: lut_13 = 8'h11;
			8'h74: lut_13 = 8'h32;
			8'h75: lut_13 = 8'h3F;
			8'h76: lut_13 = 8'h28;
			8'h77: lut_13 = 8'h25;
			8'h78: lut_13 = 8'h6E;
			8'h79: lut_13 = 8'h63;
			8'h7A: lut_13 = 8'h74;
			8'h7B: lut_13 = 8'h79;
			8'h7C: lut_13 = 8'h5A;
			8'h7D: lut_13 = 8'h57;
			8'h7E: lut_13 = 8'h40;
			8'h7F: lut_13 = 8'h4D;
			8'h80: lut_13 = 8'hDA;
			8'h81: lut_13 = 8'hD7;
			8'h82: lut_13 = 8'hC0;
			8'h83: lut_13 = 8'hCD;
			8'h84: lut_13 = 8'hEE;
			8'h85: lut_13 = 8'hE3;
			8'h86: lut_13 = 8'hF4;
			8'h87: lut_13 = 8'hF9;
			8'h88: lut_13 = 8'hB2;
			8'h89: lut_13 = 8'hBF;
			8'h8A: lut_13 = 8'hA8;
			8'h8B: lut_13 = 8'hA5;
			8'h8C: lut_13 = 8'h86;
			8'h8D: lut_13 = 8'h8B;
			8'h8E: lut_13 = 8'h9C;
			8'h8F: lut_13 = 8'h91;
			8'h90: lut_13 = 8'h0A;
			8'h91: lut_13 = 8'h07;
			8'h92: lut_13 = 8'h10;
			8'h93: lut_13 = 8'h1D;
			8'h94: lut_13 = 8'h3E;
			8'h95: lut_13 = 8'h33;
			8'h96: lut_13 = 8'h24;
			8'h97: lut_13 = 8'h29;
			8'h98: lut_13 = 8'h62;
			8'h99: lut_13 = 8'h6F;
			8'h9A: lut_13 = 8'h78;
			8'h9B: lut_13 = 8'h75;
			8'h9C: lut_13 = 8'h56;
			8'h9D: lut_13 = 8'h5B;
			8'h9E: lut_13 = 8'h4C;
			8'h9F: lut_13 = 8'h41;
			8'hA0: lut_13 = 8'h61;
			8'hA1: lut_13 = 8'h6C;
			8'hA2: lut_13 = 8'h7B;
			8'hA3: lut_13 = 8'h76;
			8'hA4: lut_13 = 8'h55;
			8'hA5: lut_13 = 8'h58;
			8'hA6: lut_13 = 8'h4F;
			8'hA7: lut_13 = 8'h42;
			8'hA8: lut_13 = 8'h09;
			8'hA9: lut_13 = 8'h04;
			8'hAA: lut_13 = 8'h13;
			8'hAB: lut_13 = 8'h1E;
			8'hAC: lut_13 = 8'h3D;
			8'hAD: lut_13 = 8'h30;
			8'hAE: lut_13 = 8'h27;
			8'hAF: lut_13 = 8'h2A;
			8'hB0: lut_13 = 8'hB1;
			8'hB1: lut_13 = 8'hBC;
			8'hB2: lut_13 = 8'hAB;
			8'hB3: lut_13 = 8'hA6;
			8'hB4: lut_13 = 8'h85;
			8'hB5: lut_13 = 8'h88;
			8'hB6: lut_13 = 8'h9F;
			8'hB7: lut_13 = 8'h92;
			8'hB8: lut_13 = 8'hD9;
			8'hB9: lut_13 = 8'hD4;
			8'hBA: lut_13 = 8'hC3;
			8'hBB: lut_13 = 8'hCE;
			8'hBC: lut_13 = 8'hED;
			8'hBD: lut_13 = 8'hE0;
			8'hBE: lut_13 = 8'hF7;
			8'hBF: lut_13 = 8'hFA;
			8'hC0: lut_13 = 8'hB7;
			8'hC1: lut_13 = 8'hBA;
			8'hC2: lut_13 = 8'hAD;
			8'hC3: lut_13 = 8'hA0;
			8'hC4: lut_13 = 8'h83;
			8'hC5: lut_13 = 8'h8E;
			8'hC6: lut_13 = 8'h99;
			8'hC7: lut_13 = 8'h94;
			8'hC8: lut_13 = 8'hDF;
			8'hC9: lut_13 = 8'hD2;
			8'hCA: lut_13 = 8'hC5;
			8'hCB: lut_13 = 8'hC8;
			8'hCC: lut_13 = 8'hEB;
			8'hCD: lut_13 = 8'hE6;
			8'hCE: lut_13 = 8'hF1;
			8'hCF: lut_13 = 8'hFC;
			8'hD0: lut_13 = 8'h67;
			8'hD1: lut_13 = 8'h6A;
			8'hD2: lut_13 = 8'h7D;
			8'hD3: lut_13 = 8'h70;
			8'hD4: lut_13 = 8'h53;
			8'hD5: lut_13 = 8'h5E;
			8'hD6: lut_13 = 8'h49;
			8'hD7: lut_13 = 8'h44;
			8'hD8: lut_13 = 8'h0F;
			8'hD9: lut_13 = 8'h02;
			8'hDA: lut_13 = 8'h15;
			8'hDB: lut_13 = 8'h18;
			8'hDC: lut_13 = 8'h3B;
			8'hDD: lut_13 = 8'h36;
			8'hDE: lut_13 = 8'h21;
			8'hDF: lut_13 = 8'h2C;
			8'hE0: lut_13 = 8'h0C;
			8'hE1: lut_13 = 8'h01;
			8'hE2: lut_13 = 8'h16;
			8'hE3: lut_13 = 8'h1B;
			8'hE4: lut_13 = 8'h38;
			8'hE5: lut_13 = 8'h35;
			8'hE6: lut_13 = 8'h22;
			8'hE7: lut_13 = 8'h2F;
			8'hE8: lut_13 = 8'h64;
			8'hE9: lut_13 = 8'h69;
			8'hEA: lut_13 = 8'h7E;
			8'hEB: lut_13 = 8'h73;
			8'hEC: lut_13 = 8'h50;
			8'hED: lut_13 = 8'h5D;
			8'hEE: lut_13 = 8'h4A;
			8'hEF: lut_13 = 8'h47;
			8'hF0: lut_13 = 8'hDC;
			8'hF1: lut_13 = 8'hD1;
			8'hF2: lut_13 = 8'hC6;
			8'hF3: lut_13 = 8'hCB;
			8'hF4: lut_13 = 8'hE8;
			8'hF5: lut_13 = 8'hE5;
			8'hF6: lut_13 = 8'hF2;
			8'hF7: lut_13 = 8'hFF;
			8'hF8: lut_13 = 8'hB4;
			8'hF9: lut_13 = 8'hB9;
			8'hFA: lut_13 = 8'hAE;
			8'hFB: lut_13 = 8'hA3;
			8'hFC: lut_13 = 8'h80;
			8'hFD: lut_13 = 8'h8D;
			8'hFE: lut_13 = 8'h9A;
			default: lut_13 = 8'h97;
		endcase
	endfunction
	
	function integer lut_14(input integer a);
		case (a)
			8'h00: lut_14 = 8'h00;
			8'h01: lut_14 = 8'h0E;
			8'h02: lut_14 = 8'h1C;
			8'h03: lut_14 = 8'h12;
			8'h04: lut_14 = 8'h38;
			8'h05: lut_14 = 8'h36;
			8'h06: lut_14 = 8'h24;
			8'h07: lut_14 = 8'h2A;
			8'h08: lut_14 = 8'h70;
			8'h09: lut_14 = 8'h7E;
			8'h0A: lut_14 = 8'h6C;
			8'h0B: lut_14 = 8'h62;
			8'h0C: lut_14 = 8'h48;
			8'h0D: lut_14 = 8'h46;
			8'h0E: lut_14 = 8'h54;
			8'h0F: lut_14 = 8'h5A;
			8'h10: lut_14 = 8'hE0;
			8'h11: lut_14 = 8'hEE;
			8'h12: lut_14 = 8'hFC;
			8'h13: lut_14 = 8'hF2;
			8'h14: lut_14 = 8'hD8;
			8'h15: lut_14 = 8'hD6;
			8'h16: lut_14 = 8'hC4;
			8'h17: lut_14 = 8'hCA;
			8'h18: lut_14 = 8'h90;
			8'h19: lut_14 = 8'h9E;
			8'h1A: lut_14 = 8'h8C;
			8'h1B: lut_14 = 8'h82;
			8'h1C: lut_14 = 8'hA8;
			8'h1D: lut_14 = 8'hA6;
			8'h1E: lut_14 = 8'hB4;
			8'h1F: lut_14 = 8'hBA;
			8'h20: lut_14 = 8'hDB;
			8'h21: lut_14 = 8'hD5;
			8'h22: lut_14 = 8'hC7;
			8'h23: lut_14 = 8'hC9;
			8'h24: lut_14 = 8'hE3;
			8'h25: lut_14 = 8'hED;
			8'h26: lut_14 = 8'hFF;
			8'h27: lut_14 = 8'hF1;
			8'h28: lut_14 = 8'hAB;
			8'h29: lut_14 = 8'hA5;
			8'h2A: lut_14 = 8'hB7;
			8'h2B: lut_14 = 8'hB9;
			8'h2C: lut_14 = 8'h93;
			8'h2D: lut_14 = 8'h9D;
			8'h2E: lut_14 = 8'h8F;
			8'h2F: lut_14 = 8'h81;
			8'h30: lut_14 = 8'h3B;
			8'h31: lut_14 = 8'h35;
			8'h32: lut_14 = 8'h27;
			8'h33: lut_14 = 8'h29;
			8'h34: lut_14 = 8'h03;
			8'h35: lut_14 = 8'h0D;
			8'h36: lut_14 = 8'h1F;
			8'h37: lut_14 = 8'h11;
			8'h38: lut_14 = 8'h4B;
			8'h39: lut_14 = 8'h45;
			8'h3A: lut_14 = 8'h57;
			8'h3B: lut_14 = 8'h59;
			8'h3C: lut_14 = 8'h73;
			8'h3D: lut_14 = 8'h7D;
			8'h3E: lut_14 = 8'h6F;
			8'h3F: lut_14 = 8'h61;
			8'h40: lut_14 = 8'hAD;
			8'h41: lut_14 = 8'hA3;
			8'h42: lut_14 = 8'hB1;
			8'h43: lut_14 = 8'hBF;
			8'h44: lut_14 = 8'h95;
			8'h45: lut_14 = 8'h9B;
			8'h46: lut_14 = 8'h89;
			8'h47: lut_14 = 8'h87;
			8'h48: lut_14 = 8'hDD;
			8'h49: lut_14 = 8'hD3;
			8'h4A: lut_14 = 8'hC1;
			8'h4B: lut_14 = 8'hCF;
			8'h4C: lut_14 = 8'hE5;
			8'h4D: lut_14 = 8'hEB;
			8'h4E: lut_14 = 8'hF9;
			8'h4F: lut_14 = 8'hF7;
			8'h50: lut_14 = 8'h4D;
			8'h51: lut_14 = 8'h43;
			8'h52: lut_14 = 8'h51;
			8'h53: lut_14 = 8'h5F;
			8'h54: lut_14 = 8'h75;
			8'h55: lut_14 = 8'h7B;
			8'h56: lut_14 = 8'h69;
			8'h57: lut_14 = 8'h67;
			8'h58: lut_14 = 8'h3D;
			8'h59: lut_14 = 8'h33;
			8'h5A: lut_14 = 8'h21;
			8'h5B: lut_14 = 8'h2F;
			8'h5C: lut_14 = 8'h05;
			8'h5D: lut_14 = 8'h0B;
			8'h5E: lut_14 = 8'h19;
			8'h5F: lut_14 = 8'h17;
			8'h60: lut_14 = 8'h76;
			8'h61: lut_14 = 8'h78;
			8'h62: lut_14 = 8'h6A;
			8'h63: lut_14 = 8'h64;
			8'h64: lut_14 = 8'h4E;
			8'h65: lut_14 = 8'h40;
			8'h66: lut_14 = 8'h52;
			8'h67: lut_14 = 8'h5C;
			8'h68: lut_14 = 8'h06;
			8'h69: lut_14 = 8'h08;
			8'h6A: lut_14 = 8'h1A;
			8'h6B: lut_14 = 8'h14;
			8'h6C: lut_14 = 8'h3E;
			8'h6D: lut_14 = 8'h30;
			8'h6E: lut_14 = 8'h22;
			8'h6F: lut_14 = 8'h2C;
			8'h70: lut_14 = 8'h96;
			8'h71: lut_14 = 8'h98;
			8'h72: lut_14 = 8'h8A;
			8'h73: lut_14 = 8'h84;
			8'h74: lut_14 = 8'hAE;
			8'h75: lut_14 = 8'hA0;
			8'h76: lut_14 = 8'hB2;
			8'h77: lut_14 = 8'hBC;
			8'h78: lut_14 = 8'hE6;
			8'h79: lut_14 = 8'hE8;
			8'h7A: lut_14 = 8'hFA;
			8'h7B: lut_14 = 8'hF4;
			8'h7C: lut_14 = 8'hDE;
			8'h7D: lut_14 = 8'hD0;
			8'h7E: lut_14 = 8'hC2;
			8'h7F: lut_14 = 8'hCC;
			8'h80: lut_14 = 8'h41;
			8'h81: lut_14 = 8'h4F;
			8'h82: lut_14 = 8'h5D;
			8'h83: lut_14 = 8'h53;
			8'h84: lut_14 = 8'h79;
			8'h85: lut_14 = 8'h77;
			8'h86: lut_14 = 8'h65;
			8'h87: lut_14 = 8'h6B;
			8'h88: lut_14 = 8'h31;
			8'h89: lut_14 = 8'h3F;
			8'h8A: lut_14 = 8'h2D;
			8'h8B: lut_14 = 8'h23;
			8'h8C: lut_14 = 8'h09;
			8'h8D: lut_14 = 8'h07;
			8'h8E: lut_14 = 8'h15;
			8'h8F: lut_14 = 8'h1B;
			8'h90: lut_14 = 8'hA1;
			8'h91: lut_14 = 8'hAF;
			8'h92: lut_14 = 8'hBD;
			8'h93: lut_14 = 8'hB3;
			8'h94: lut_14 = 8'h99;
			8'h95: lut_14 = 8'h97;
			8'h96: lut_14 = 8'h85;
			8'h97: lut_14 = 8'h8B;
			8'h98: lut_14 = 8'hD1;
			8'h99: lut_14 = 8'hDF;
			8'h9A: lut_14 = 8'hCD;
			8'h9B: lut_14 = 8'hC3;
			8'h9C: lut_14 = 8'hE9;
			8'h9D: lut_14 = 8'hE7;
			8'h9E: lut_14 = 8'hF5;
			8'h9F: lut_14 = 8'hFB;
			8'hA0: lut_14 = 8'h9A;
			8'hA1: lut_14 = 8'h94;
			8'hA2: lut_14 = 8'h86;
			8'hA3: lut_14 = 8'h88;
			8'hA4: lut_14 = 8'hA2;
			8'hA5: lut_14 = 8'hAC;
			8'hA6: lut_14 = 8'hBE;
			8'hA7: lut_14 = 8'hB0;
			8'hA8: lut_14 = 8'hEA;
			8'hA9: lut_14 = 8'hE4;
			8'hAA: lut_14 = 8'hF6;
			8'hAB: lut_14 = 8'hF8;
			8'hAC: lut_14 = 8'hD2;
			8'hAD: lut_14 = 8'hDC;
			8'hAE: lut_14 = 8'hCE;
			8'hAF: lut_14 = 8'hC0;
			8'hB0: lut_14 = 8'h7A;
			8'hB1: lut_14 = 8'h74;
			8'hB2: lut_14 = 8'h66;
			8'hB3: lut_14 = 8'h68;
			8'hB4: lut_14 = 8'h42;
			8'hB5: lut_14 = 8'h4C;
			8'hB6: lut_14 = 8'h5E;
			8'hB7: lut_14 = 8'h50;
			8'hB8: lut_14 = 8'h0A;
			8'hB9: lut_14 = 8'h04;
			8'hBA: lut_14 = 8'h16;
			8'hBB: lut_14 = 8'h18;
			8'hBC: lut_14 = 8'h32;
			8'hBD: lut_14 = 8'h3C;
			8'hBE: lut_14 = 8'h2E;
			8'hBF: lut_14 = 8'h20;
			8'hC0: lut_14 = 8'hEC;
			8'hC1: lut_14 = 8'hE2;
			8'hC2: lut_14 = 8'hF0;
			8'hC3: lut_14 = 8'hFE;
			8'hC4: lut_14 = 8'hD4;
			8'hC5: lut_14 = 8'hDA;
			8'hC6: lut_14 = 8'hC8;
			8'hC7: lut_14 = 8'hC6;
			8'hC8: lut_14 = 8'h9C;
			8'hC9: lut_14 = 8'h92;
			8'hCA: lut_14 = 8'h80;
			8'hCB: lut_14 = 8'h8E;
			8'hCC: lut_14 = 8'hA4;
			8'hCD: lut_14 = 8'hAA;
			8'hCE: lut_14 = 8'hB8;
			8'hCF: lut_14 = 8'hB6;
			8'hD0: lut_14 = 8'h0C;
			8'hD1: lut_14 = 8'h02;
			8'hD2: lut_14 = 8'h10;
			8'hD3: lut_14 = 8'h1E;
			8'hD4: lut_14 = 8'h34;
			8'hD5: lut_14 = 8'h3A;
			8'hD6: lut_14 = 8'h28;
			8'hD7: lut_14 = 8'h26;
			8'hD8: lut_14 = 8'h7C;
			8'hD9: lut_14 = 8'h72;
			8'hDA: lut_14 = 8'h60;
			8'hDB: lut_14 = 8'h6E;
			8'hDC: lut_14 = 8'h44;
			8'hDD: lut_14 = 8'h4A;
			8'hDE: lut_14 = 8'h58;
			8'hDF: lut_14 = 8'h56;
			8'hE0: lut_14 = 8'h37;
			8'hE1: lut_14 = 8'h39;
			8'hE2: lut_14 = 8'h2B;
			8'hE3: lut_14 = 8'h25;
			8'hE4: lut_14 = 8'h0F;
			8'hE5: lut_14 = 8'h01;
			8'hE6: lut_14 = 8'h13;
			8'hE7: lut_14 = 8'h1D;
			8'hE8: lut_14 = 8'h47;
			8'hE9: lut_14 = 8'h49;
			8'hEA: lut_14 = 8'h5B;
			8'hEB: lut_14 = 8'h55;
			8'hEC: lut_14 = 8'h7F;
			8'hED: lut_14 = 8'h71;
			8'hEE: lut_14 = 8'h63;
			8'hEF: lut_14 = 8'h6D;
			8'hF0: lut_14 = 8'hD7;
			8'hF1: lut_14 = 8'hD9;
			8'hF2: lut_14 = 8'hCB;
			8'hF3: lut_14 = 8'hC5;
			8'hF4: lut_14 = 8'hEF;
			8'hF5: lut_14 = 8'hE1;
			8'hF6: lut_14 = 8'hF3;
			8'hF7: lut_14 = 8'hFD;
			8'hF8: lut_14 = 8'hA7;
			8'hF9: lut_14 = 8'hA9;
			8'hFA: lut_14 = 8'hBB;
			8'hFB: lut_14 = 8'hB5;
			8'hFC: lut_14 = 8'h9F;
			8'hFD: lut_14 = 8'h91;
			8'hFE: lut_14 = 8'h83;
			default: lut_14 = 8'h8D;
		endcase

	endfunction
endmodule
